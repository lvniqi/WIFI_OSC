library verilog;
use verilog.vl_types.all;
entity fifo_control is
    port(
        clk             : in     vl_logic
    );
end fifo_control;
